@00000000
0F 00 0F 00 0F 00 01 20 00 00 00 01 01 30 00 00 
00 02 0E 22 C0 03 03 00 00 00 19 B6 0E 23 C0 03 
1A 00 00 00 10 2C 03 00 00 00 19 B6 0E 23 C4 03 
03 00 00 00 19 B6 0E 22 C4 03 1A 00 00 00 10 46 
03 00 00 00 19 B6 01 20 A0 00 01 00 01 30 A0 00 
02 00 0E 32 D4 03 03 00 00 00 19 B6 0E 23 D4 03 
1A 00 00 00 10 6C 03 00 00 00 19 B6 0E 22 D4 03 
1A 00 00 00 10 7C 03 00 00 00 19 B6 0E 23 D0 03 
03 00 00 00 19 B6 0E 32 D0 03 1A 00 00 00 10 96 
03 00 00 00 19 B6 0E 22 D0 03 1A 00 00 00 10 A6 
03 00 00 00 19 B6 0E 32 E0 03 03 00 00 00 19 B6 
0E 23 E0 03 1A 00 00 00 10 C0 03 00 00 00 19 B6 
0E 22 E0 03 03 00 00 00 19 B6 0E 23 E4 03 03 00 
00 00 19 B6 0E 32 E4 03 1A 00 00 00 10 E4 03 00 
00 00 19 B6 0E 22 E4 03 03 00 00 00 19 B6 01 20 
FF FF FF 9C 01 30 00 00 00 64 0E 32 CC 03 03 00 
00 00 19 B6 0E 23 CC 03 1A 00 00 00 11 14 03 00 
00 00 19 B6 0E 22 CC 03 1A 00 00 00 11 24 03 00 
00 00 19 B6 0E 23 C8 03 03 00 00 00 19 B6 0E 32 
C8 03 1A 00 00 00 11 3E 03 00 00 00 19 B6 0E 22 
C8 03 1A 00 00 00 11 4E 03 00 00 00 19 B6 0E 32 
D8 03 03 00 00 00 19 B6 0E 23 D8 03 1A 00 00 00 
11 68 03 00 00 00 19 B6 0E 22 D8 03 03 00 00 00 
19 B6 0E 23 DC 03 03 00 00 00 19 B6 0E 32 DC 03 
1A 00 00 00 11 8C 03 00 00 00 19 B6 0E 22 DC 03 
03 00 00 00 19 B6 01 20 00 00 00 00 01 30 00 00 
00 C8 01 40 00 00 00 C8 02 23 0E 24 C0 03 03 00 
00 00 19 B6 01 20 00 00 00 64 01 30 00 00 00 C8 
01 40 00 00 01 2C 05 23 0E 24 C0 03 03 00 00 00 
19 B6 01 20 00 00 01 2C 01 30 00 00 00 64 01 40 
00 00 00 C8 29 23 0E 24 C0 03 03 00 00 00 19 B6 
01 20 12 34 56 78 01 30 F0 F0 F0 F0 01 40 10 30 
50 70 26 23 0E 24 C0 03 03 00 00 00 19 B6 01 20 
12 34 01 01 01 30 FF F0 10 10 01 40 FF F4 11 11 
2B 23 0E 24 C0 03 03 00 00 00 19 B6 01 20 12 34 
01 01 01 30 FF F0 10 10 01 40 ED C4 11 11 2E 23 
0E 24 C0 03 03 00 00 00 19 B6 01 20 00 00 00 00 
01 30 12 34 56 78 01 40 ED CB A9 87 2C 23 0E 24 
C0 03 03 00 00 00 19 B6 01 20 00 00 00 00 01 30 
00 00 00 64 01 40 FF FF FF 9C 2A 23 0E 24 C0 03 
03 00 00 00 19 B6 01 20 00 00 00 00 01 30 FF FF 
FF 9C 01 40 00 00 00 64 2A 23 0E 24 C0 03 03 00 
00 00 19 B6 01 20 00 00 00 64 01 40 00 00 01 5E 
82 FA 0E 24 C0 03 03 00 00 00 19 B6 01 20 00 00 
01 90 01 40 00 00 00 96 92 FA 0E 24 C0 03 03 00 
00 00 19 B6 01 20 00 AA AA 00 01 30 00 00 00 05 
01 40 00 05 55 50 27 23 0E 24 C0 03 03 00 00 00 
19 B6 01 20 00 55 55 00 01 30 00 00 00 05 01 40 
0A AA A0 00 28 23 0E 24 C0 03 03 00 00 00 19 B6 
01 20 00 AA AA 00 01 30 00 00 00 05 01 40 00 05 
55 50 2D 23 0E 24 C0 03 03 00 00 00 19 B6 01 20 
80 AA AA 00 01 30 00 00 00 05 01 40 FC 05 55 50 
2D 23 0E 24 C0 03 03 00 00 00 19 B6 01 20 00 00 
00 64 01 30 00 00 00 C8 01 40 00 00 4E 20 2F 23 
0E 24 C0 03 03 00 00 00 19 B6 01 20 00 00 00 64 
01 30 FF FF FF 38 01 40 FF FF B1 E0 2F 23 0E 24 
C0 03 03 00 00 00 19 B6 01 20 FF FF FF 9C 01 30 
00 00 00 C8 01 40 FF FF B1 E0 2F 23 0E 24 C0 03 
03 00 00 00 19 B6 01 20 FF FF FF 9C 01 30 FF FF 
FF 38 01 40 00 00 4E 20 2F 23 0E 24 C0 03 03 00 
00 00 19 B6 01 20 00 00 4E 20 01 30 00 00 00 C8 
01 40 00 00 00 64 31 23 0E 24 C0 03 03 00 00 00 
19 B6 01 20 00 00 4E 20 01 30 FF FF FF 38 01 40 
FF FF FF 9C 31 23 0E 24 C0 03 03 00 00 00 19 B6 
01 20 FF FF B1 E0 01 30 00 00 00 C8 01 40 FF FF 
FF 9C 31 23 0E 24 C0 03 03 00 00 00 19 B6 01 20 
FF FF B1 E0 01 30 FF FF FF 38 01 40 00 00 00 64 
31 23 0E 24 C0 03 03 00 00 00 19 B6 01 20 B2 D0 
5E 00 01 30 08 F0 D1 80 01 40 00 00 00 14 32 23 
0E 24 C0 03 03 00 00 00 19 B6 01 20 00 00 4E 2A 
01 30 00 00 00 C8 01 40 00 00 00 0A 33 23 0E 24 
C0 03 03 00 00 00 19 B6 01 20 00 00 4E 2A 01 30 
FF FF FF 38 01 40 00 00 00 0A 33 23 0E 24 C0 03 
03 00 00 00 19 B6 01 20 FF FF B1 D6 01 30 00 00 
00 C8 01 40 FF FF FF F6 33 23 0E 24 C0 03 03 00 
00 00 19 B6 01 20 FF FF B1 D6 01 30 FF FF FF 38 
01 40 FF FF FF F6 33 23 0E 24 C0 03 03 00 00 00 
19 B6 01 20 B2 D0 5E 64 01 30 08 F0 D1 80 01 40 
00 00 00 64 34 23 0E 24 C0 03 03 00 00 00 19 B6 
01 30 12 34 56 78 09 30 00 20 0A 00 08 40 00 20 
0A 00 0E 34 C0 03 03 00 00 00 19 B6 2E 44 22 40 
00 20 0A 00 01 50 00 00 12 34 0E 45 C0 03 03 00 
00 00 19 B6 2E 44 22 40 00 20 0A 02 01 50 00 00 
56 78 0E 45 C0 03 03 00 00 00 19 B6 1D 40 00 20 
0A 00 01 50 00 00 00 12 0E 45 C0 03 03 00 00 00 
19 B6 1D 40 00 20 0A 01 01 50 00 00 00 34 0E 45 
C0 03 03 00 00 00 19 B6 1D 40 00 20 0A 02 01 50 
00 00 00 56 0E 45 C0 03 03 00 00 00 19 B6 1D 40 
00 20 0A 03 01 50 00 00 00 78 0E 45 C0 03 03 00 
00 00 19 B6 01 30 12 34 56 78 09 30 00 20 0A 01 
08 40 00 20 0A 01 0E 34 C0 03 03 00 00 00 19 B6 
2E 44 22 40 00 20 0A 01 01 50 00 00 12 34 0E 45 
C0 03 03 00 00 00 19 B6 2E 44 22 40 00 20 0A 03 
01 50 00 00 56 78 0E 45 C0 03 03 00 00 00 19 B6 
1D 40 00 20 0A 01 01 50 00 00 00 12 0E 45 C0 03 
03 00 00 00 19 B6 1D 40 00 20 0A 02 01 50 00 00 
00 34 0E 45 C0 03 03 00 00 00 19 B6 1D 40 00 20 
0A 03 01 50 00 00 00 56 0E 45 C0 03 03 00 00 00 
19 B6 1D 40 00 20 0A 04 01 50 00 00 00 78 0E 45 
C0 03 03 00 00 00 19 B6 01 30 00 00 12 34 24 30 
00 20 0A 00 22 40 00 20 0A 00 0E 34 C0 03 03 00 
00 00 19 B6 1D 40 00 20 0A 00 01 50 00 00 00 12 
0E 45 C0 03 03 00 00 00 19 B6 1D 40 00 20 0A 01 
01 50 00 00 00 34 0E 45 C0 03 03 00 00 00 19 B6 
01 30 00 00 12 34 24 30 00 20 0A 01 22 40 00 20 
0A 01 0E 34 C0 03 03 00 00 00 19 B6 1D 40 00 20 
0A 01 01 50 00 00 00 12 0E 45 C0 03 03 00 00 00 
19 B6 1D 40 00 20 0A 02 01 50 00 00 00 34 0E 45 
C0 03 03 00 00 00 19 B6 01 30 00 00 00 12 1F 30 
00 20 0A 00 1D 40 00 20 0A 00 0E 34 C0 03 03 00 
00 00 19 B6 01 30 00 00 00 12 1F 30 00 20 0A 01 
1D 40 00 20 0A 01 0E 34 C0 03 03 00 00 00 19 B6 
01 30 AA AA AA AA 09 30 00 20 0A 00 09 30 00 20 
0A 04 01 30 12 34 56 78 09 30 00 20 0A 01 1D 30 
00 20 0A 00 01 40 00 00 00 AA 0E 34 C0 03 03 00 
00 00 19 B6 1D 30 00 20 0A 05 0E 34 C0 03 03 00 
00 00 19 B6 01 30 AA AA AA AA 09 30 00 20 0A 00 
01 30 00 00 12 34 24 30 00 20 0A 01 1D 30 00 20 
0A 00 01 40 00 00 00 AA 0E 34 C0 03 03 00 00 00 
19 B6 1D 30 00 20 0A 03 0E 34 C0 03 03 00 00 00 
19 B6 01 30 AA AA AA AA 09 30 00 20 0A 00 01 30 
00 00 00 12 1F 30 00 20 0A 00 1D 30 00 20 0A 01 
01 40 00 00 00 AA 0E 34 C0 03 03 00 00 00 19 B6 
01 30 AA AA AA AA 09 30 00 20 0A 00 01 30 00 00 
00 12 1F 30 00 20 0A 01 1D 30 00 20 0A 00 01 40 
00 00 00 AA 0E 34 C0 03 03 00 00 00 19 B6 01 30 
00 20 0A 10 01 40 12 34 56 78 0B 34 0A 53 0E 54 
C0 03 03 00 00 00 19 B6 08 50 00 20 0A 10 0E 54 
C0 03 03 00 00 00 19 B6 01 30 00 20 0A 20 01 40 
00 00 12 34 23 34 21 53 0E 54 C0 03 03 00 00 00 
19 B6 22 50 00 20 0A 20 0E 54 C0 03 03 00 00 00 
19 B6 01 30 00 20 0A 30 01 40 00 00 00 12 1E 34 
1C 53 0E 54 C0 03 03 00 00 00 19 B6 1D 50 00 20 
0A 30 0E 54 C0 03 03 00 00 00 19 B6 01 30 00 20 
0B 10 01 40 12 34 56 78 0D 34 00 00 01 00 0C 53 
00 00 01 00 0E 54 C0 03 03 00 00 00 19 B6 08 50 
00 20 0C 10 0E 54 C0 03 03 00 00 00 19 B6 01 30 
00 20 0B 20 01 40 00 00 12 34 39 34 00 00 01 00 
38 53 00 00 01 00 0E 54 C0 03 03 00 00 00 19 B6 
22 50 00 20 0C 20 0E 54 C0 03 03 00 00 00 19 B6 
01 30 00 20 0B 30 01 40 00 00 00 12 37 34 00 00 
01 00 36 53 00 00 01 00 0E 54 C0 03 03 00 00 00 
19 B6 1D 50 00 20 0C 30 0E 54 C0 03 03 00 00 00 
19 B6 01 20 00 00 09 00 25 20 03 00 00 00 19 B6 
1A 00 00 00 19 0C 03 00 00 00 19 B6 01 10 00 20 
0A 80 01 30 00 00 00 64 06 13 01 50 00 20 0A 7C 
0E 15 C0 03 03 00 00 00 19 B6 07 14 0E 34 C0 03 
03 00 00 00 19 B6 01 50 00 20 0A 80 0E 15 C0 03 
03 00 00 00 19 B6 1A 00 00 00 19 64 06 12 0C 30 
00 00 00 0C 0C 40 00 00 00 10 05 34 02 E0 9E 04 
07 E2 04 00 01 30 00 00 03 E8 06 13 01 30 00 00 
01 F4 06 13 03 00 00 00 19 4C 01 40 00 00 05 DC 
0E 34 C0 03 03 00 00 00 19 B6 01 30 00 00 07 D0 
06 13 01 30 00 00 03 E8 06 13 01 30 00 00 09 4C 
19 30 01 40 00 00 0B B8 0E 34 C0 03 03 00 00 00 
19 B6 2E 22 04 00 0C 21 00 00 00 04 80 0C 04 00 
