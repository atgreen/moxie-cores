@30000000
01 10 30 FF 8C 54 2E 00 01 20 30 00 0B CC 01 30
30 00 0C 54 2E 44 0E 23 C0 06 0D 24 00 00 82 04
1A 00 30 00 00 16 01 20 00 00 FE ED 24 20 F0 00
00 00 2E 22 2E 33 2E 44 03 00 30 00 06 64 1A 00
30 00 00 3E 01 30 00 00 00 01 22 20 F0 00 00 08
0E 23 C7 FB 22 20 F0 00 00 0C 04 00 6D 6F 78 69
65 00 91 18 01 30 30 00 0B C8 01 20 30 00 0B C8
0E 32 C0 07 01 30 00 00 00 00 2E 44 0E 34 C0 01
19 30 04 00 91 18 01 40 30 00 0B C8 01 20 30 00
0B C8 29 42 01 30 00 00 00 02 2D 43 01 50 00 00
00 1F 02 34 27 35 05 34 01 40 00 00 00 01 2D 34
2E 55 0E 35 C0 06 01 40 00 00 00 00 0E 45 C0 01
19 40 04 00 06 18 06 19 06 1A 91 18 1D 30 30 00
0B CC 2E 22 0E 32 C4 33 01 A0 00 00 00 02 01 80
30 00 0B C0 01 20 30 00 0B BC 29 82 2D 8A 98 01
02 92 08 20 30 00 0B D0 0E 28 E0 0E 82 01 09 20
30 00 0B D0 28 2A 02 39 05 32 0A 23 19 20 08 20
30 00 0B D0 0E 28 D3 F2 03 00 30 00 00 62 01 30
00 00 00 00 2E 22 0E 32 C0 04 01 20 30 00 0B C4
19 30 1B 20 00 00 00 01 1F 20 30 00 0B CC 02 E0
9E 0C 07 EA 07 E9 07 E8 04 00 91 18 04 00 91 18
01 40 00 00 00 00 2E 22 0E 42 C0 07 01 30 30 00
0B D4 01 20 30 00 0B C4 19 40 03 00 30 00 00 84
04 00 91 18 04 00 06 18 2E 88 01 60 F0 00 00 08
01 E0 00 00 00 01 1C 42 0E 48 C4 04 02 E0 9E 04
07 E8 04 00 38 56 00 02 11 55 0E 5E C7 FB 39 64
00 06 0E 3E C4 07 08 50 30 00 0C 4C 05 54 09 50
30 00 0C 4C 82 01 1A 00 30 00 01 86 02 32 12 22
01 40 00 00 00 46 0E 24 D4 10 01 40 00 00 00 40
0E 24 D4 16 93 30 12 33 01 40 00 00 00 09 0E 34
E4 0D 01 20 FF FF FF FF 04 00 93 61 12 33 01 40
00 00 00 05 0E 34 D7 F5 92 57 04 00 92 30 04 00
92 37 04 00 06 18 06 19 06 1A 91 18 02 92 2E 88
01 A0 FF FF FF FF 99 01 0E 9A C4 07 02 28 02 E0
9E 0C 07 EA 07 E9 07 E8 04 00 03 00 30 00 00 44
12 22 03 00 30 00 01 BC 01 30 00 00 00 04 28 83
05 82 1A 00 30 00 02 16 06 18 06 19 91 18 2E 88
01 90 30 00 00 44 19 90 12 22 03 00 30 00 01 BC
2E 33 0E 23 C8 08 01 30 00 00 00 04 28 83 05 82
1A 00 30 00 02 56 02 28 02 E0 9E 08 07 E9 07 E8
04 00 06 18 06 19 06 1A 01 40 30 00 0B EC 01 30
00 00 00 1C 02 64 01 A0 00 00 00 0F 01 90 30 00
0A C0 01 E0 FF FF FF FC 02 52 2D 53 26 5A 02 89
05 85 1C 58 1E 45 93 04 84 01 0E 3E C7 F5 2E 22
37 62 00 08 01 20 30 00 0B EC 02 E0 9E 0C 07 EA
07 E9 07 E8 04 00 02 32 01 20 30 00 0B F8 01 40
00 00 00 04 02 53 2D 54 01 60 00 00 00 0F 26 56
01 40 30 00 0A C0 02 E4 05 E5 1C 5E 1E 25 26 36
05 43 1C 34 37 23 00 01 2E 33 37 23 00 02 04 00
06 18 91 18 01 80 30 00 01 76 2E 33 01 20 30 00
0A D4 19 80 08 20 30 00 0C 4C 03 00 30 00 02 D6
2E 33 19 80 2E 22 09 20 30 00 0C 4C 02 E0 9E 04
07 E8 04 00 06 18 06 19 06 1A 06 1B 06 1C 91 18
2E 88 22 30 30 00 0C 50 11 23 0E 28 01 90 30 00
00 44 C4 31 01 A0 00 00 00 24 19 90 12 22 0E 2A
C7 FC 19 90 12 22 01 30 00 00 00 63 0E 23 C0 5A
D4 28 01 30 00 00 00 4D 0E 23 C0 AA 01 30 00 00
00 50 0E 23 C0 CD 01 30 00 00 00 3F 0E 23 C0 DC
01 A0 00 00 00 23 19 90 12 22 0E 2A C7 FC 19 90
19 90 02 38 01 20 30 00 0A E8 03 00 30 00 01 76
1A 00 30 00 03 52 24 80 30 00 0C 50 1A 00 30 00
03 72 01 30 00 00 00 6D 0E 23 C0 5D 01 30 00 00
00 70 0E 23 C0 36 01 30 00 00 00 67 0E 23 C7 D8
19 90 19 90 19 90 01 A0 30 00 01 76 02 38 01 20
30 00 0A DC 19 A0 01 90 30 00 0B FC 02 B9 8B 48
01 C0 30 00 02 82 0A 29 19 C0 01 30 00 00 00 01
19 A0 89 04 0E 9B C7 F7 03 00 30 00 03 10 1A 00
30 00 03 52 2E 33 01 20 30 00 0A D8 03 00 30 00
01 76 02 E0 9E 14 07 EC 07 EB 07 EA 07 E9 07 E8
04 00 03 00 30 00 02 48 02 A2 19 90 19 90 01 90
30 00 01 76 02 38 01 20 30 00 0A DC 19 90 01 30
00 00 00 02 02 2A 28 23 01 30 30 00 0B FC 05 32
0A 23 03 00 30 00 02 82 01 30 00 00 00 01 19 90
1A 00 30 00 04 28 01 A0 30 00 02 48 19 A0 02 B2
19 A0 02 A2 19 90 19 90 01 90 30 00 01 76 02 38
01 20 30 00 0A DC 19 90 02 CB 05 CA 02 2C 29 2B
0E 28 DF B2 02 AB 8A 01 1C 2B 03 00 30 00 02 D6
01 30 00 00 00 01 19 90 02 BA 1A 00 30 00 04 BC
01 90 30 00 02 48 19 90 02 A2 19 90 02 9A 05 92
02 29 29 2A 0E 28 CC 11 01 90 30 00 01 76 02 38
01 20 30 00 0A DC 19 90 01 30 00 00 00 01 01 20
30 00 0A E0 1A 00 30 00 04 8E 01 20 00 00 00 02
03 00 30 00 02 04 1E A2 8A 01 1A 00 30 00 04 F0
01 A0 30 00 02 48 19 A0 02 B2 19 A0 01 30 00 00
00 02 28 B3 01 30 30 00 0B FC 05 3B 0B 32 19 90
19 90 1A 00 30 00 04 F8 19 90 19 90 19 90 01 90
30 00 01 76 02 38 01 20 30 00 0A DC 19 90 01 30
00 00 00 01 01 20 30 00 0A E4 1A 00 30 00 04 8E
06 18 06 19 06 1A 06 1B 06 1C 91 18 02 82 01 20
00 00 00 04 0E 32 CC 10 01 20 00 00 00 02 0E 32
CC 04 C0 18 2E 22 0E 32 C8 0C 2E 22 24 20 F0 00
00 00 1A 00 30 00 05 B2 01 20 00 00 00 05 0E 32
C0 16 20 20 FF FF FF FF 24 20 F0 00 00 00 1A 00
30 00 05 CE 2E 22 24 20 F0 00 00 10 02 28 02 E0
9E 14 07 EC 07 EB 07 EA 07 E9 07 E8 04 00 02 A0
01 90 30 00 01 76 2E 33 01 20 30 00 0A F0 19 90
01 30 00 00 00 01 01 20 30 00 0A E4 19 90 03 00
30 00 03 10 02 9A 89 0C 01 B0 30 00 0C 04 02 CA
8C 44 02 3B 02 29 0A 42 0B 34 82 04 83 04 0E 2C
C7 FA 0A 2A 01 A0 30 00 0B FC 0D A2 00 04 0A 22
0B A2 98 02 0D A8 00 40 03 00 30 00 03 44 0A 2B
0B 92 8B 04 89 04 0E 9C C7 FA 0C 8A 00 40 1A 00
30 00 05 DC 06 18 06 19 06 1A 06 1B 06 1C 06 1D
91 24 01 C0 F0 00 00 08 20 20 00 00 00 58 39 C2
00 06 20 20 00 00 00 59 39 C2 00 06 20 20 00 00
00 5A 39 C2 00 06 01 20 30 00 08 F4 B2 01 01 90
00 00 00 01 B9 00 2E 88 09 80 30 00 0C 4C 01 A0
30 00 01 76 02 38 01 20 30 00 0A F4 19 A0 02 38
01 20 30 00 0B 14 19 A0 02 38 01 20 30 00 0B 8C
19 A0 02 38 01 20 30 00 0B 50 19 A0 24 90 30 00
0C 50 01 D0 30 00 00 44 19 D0 12 22 01 30 00 00
00 24 0E 23 C0 E8 01 30 00 00 00 53 0E 23 C7 F4
20 90 00 00 00 01 2E BB 22 30 30 00 0C 50 11 23
0E 2B C4 1D 01 80 00 00 00 53 19 D0 12 22 0E 28
C7 FC 19 D0 12 A2 02 3A 02 2A 92 30 13 22 01 50
00 00 00 09 0E 25 E4 11 01 20 00 00 00 08 28 32
05 39 24 30 F0 00 00 00 1A 00 30 00 07 48 24 B0
30 00 0C 50 1A 00 30 00 07 22 01 80 30 00 02 04
01 20 00 00 00 02 0D 03 FF E0 19 80 02 52 24 90
F0 00 00 00 01 20 00 00 00 37 0E A2 0C 30 FF E0
C0 8A D4 15 01 20 00 00 00 30 0E A2 C0 2C 01 20
00 00 00 33 0E A2 C0 39 01 20 00 00 00 08 28 32
05 39 24 30 F0 00 00 00 1A 00 30 00 07 A8 01 20
00 00 00 39 0E A2 C7 F0 2E 33 21 2C 11 22 0E 23
C4 7B 01 20 30 00 0B 90 03 00 30 00 01 76 20 20
00 00 30 00 24 20 F0 00 00 00 1A 00 30 00 00 00
1A 00 30 00 07 E0 02 25 05 25 02 82 13 28 0E 2B
C4 07 02 2B 89 01 0E 2B C3 87 1A 00 30 00 07 B8
19 D0 98 01 1A 00 30 00 07 EC 01 20 00 00 00 08
0D 05 FF DC 19 80 02 A2 0C 50 FF DC 95 04 01 30
00 00 00 04 11 25 0E 23 CC 12 01 30 00 00 00 02
11 25 0E 23 CC 1E C4 03 02 23 19 80 1E A2 01 20
00 00 00 02 19 80 89 01 1A 00 30 00 07 08 01 20
00 00 00 08 0D 03 FF E0 0D 05 FF DC 19 80 0B A2
8A 04 0C 50 FF DC 95 04 0C 30 FF E0 1A 00 30 00
08 24 01 20 00 00 00 04 0D 03 FF E0 0D 05 FF DC
19 80 23 A2 8A 02 0C 50 FF DC 95 02 0C 30 FF E0
1A 00 30 00 08 30 02 25 05 25 02 82 13 28 0E 2B
C4 06 01 20 00 00 00 01 1A 00 30 00 07 F4 19 D0
98 01 1A 00 30 00 08 9C 38 2C 00 04 39 02 FF E6
1A 00 30 00 07 BA 20 20 FF FF DE B2 24 20 F0 00
00 00 01 80 30 00 0B FC 01 40 00 00 00 50 2E 33
02 28 03 00 30 00 09 56 03 00 30 00 03 44 0C 88
00 40 25 80 91 0C 0B 10 02 01 06 1F 06 1E 06 1D
06 1C 06 1B 06 1A 06 19 06 18 06 17 06 16 06 15
06 14 06 13 06 12 A2 05 A3 02 A4 03 03 00 30 00
05 80 0D 02 00 04 01 60 00 00 00 01 A5 00 2B 56
B5 00 02 20 92 38 02 12 07 12 07 13 07 14 07 15
07 16 07 17 07 18 07 19 07 1A 07 1B 07 1C 07 1D
07 1E 07 1F 04 00 06 18 06 19 06 1A 06 1B 02 E2
01 90 00 00 00 03 02 52 26 59 2E 88 0E 58 C0 7D
02 64 96 01 0E 48 C0 6B 02 A3 02 52 01 B0 FF FF
FF FF 1A 00 30 00 09 90 96 01 8E 01 0E 6B C0 5F
85 01 1E EA 02 45 26 49 0E 48 C7 F6 01 40 00 00
00 03 0E 64 E4 4B 12 83 01 90 00 00 00 08 02 48
28 49 2B 48 01 90 00 00 00 10 02 84 28 89 2B 84
01 40 00 00 00 0F 02 A6 0E 64 E4 21 9A 10 01 40
00 00 00 04 27 A4 8A 01 28 A4 2E 99 02 45 05 49
0B 48 0D 48 00 04 0D 48 00 08 0D 48 00 0C 89 10
0E 9A C7 F4 05 59 01 40 00 00 00 0F 02 A6 26 A4
01 40 00 00 00 0C 26 64 2E 44 0E 64 C0 27 02 45
02 B5 05 BA 01 90 00 00 00 03 0B 48 84 04 02 6B
29 64 0E 69 D7 FA 02 4A 94 04 01 60 00 00 00 02
27 46 84 01 28 46 05 54 02 6A 26 69 2E 44 0E 64
C0 06 02 45 05 46 1E 53 85 01 0E 45 C7 FC 02 E0
9E 10 07 EB 07 EA 07 E9 07 E8 04 00 02 6A 2E 44
0E 64 C7 EF 1A 00 30 00 0A 4E 02 52 02 64 1A 00
30 00 09 9C 06 18 06 19 91 18 01 80 30 00 0B B8
0C 28 FF FC 01 90 FF FF FF FF 0E 29 C0 06 98 04
19 20 98 04 0A 28 0E 29 C7 FB 02 E0 9E 08 07 E9
07 E8 04 00 91 18 04 00 03 00 30 00 01 4E 03 00
30 00 0A 74 04 00 03 00 30 00 00 C4 04 00 00 00
@30000AC0
30 31 32 33 34 35 36 37 38 39 41 42 43 44 45 46
00 00 00 00 23 00 00 00 2B 00 00 00 2B 24 00 00
4F 4B 00 00 53 30 35 00 2B 24 23 30 30 00 00 00
24 00 00 00 4D 4F 58 49 45 20 4F 6E 2D 43 68 69
70 20 42 6F 6F 74 6C 6F 61 64 65 72 20 76 32 2E
30 0A 0D 00 43 6F 70 79 72 69 67 68 74 20 28 63
29 20 32 30 31 33 20 41 6E 74 68 6F 6E 79 20 47
72 65 65 6E 20 3C 67 72 65 65 6E 40 6D 6F 78 69
65 6C 6F 67 69 63 2E 63 6F 6D 3E 0A 0D 00 00 00
57 61 69 74 69 6E 67 20 66 6F 72 20 61 6E 20 53
2D 52 65 63 6F 72 64 20 44 6F 77 6E 6C 6F 61 64
20 6F 72 20 52 65 6D 6F 74 65 20 47 44 42 20 43
6F 6E 6E 65 63 74 69 6F 6E 2E 2E 2E 0A 0D 00 00
4A 75 6D 70 69 6E 67 20 74 6F 20 63 6F 64 65 20
61 74 20 30 78 33 30 30 30 30 30 30 30 2E 0A 0D
00 00 00 00 FF FF FF FF 00 00 00 00 FF FF FF FF
00 00 00 00 00 00 00 00
@30000BC8
00 00 00 00
