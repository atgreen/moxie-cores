@00000000
2B 3B 24 23 30 30 3B 24 53 30 30 23 42 33 3B
