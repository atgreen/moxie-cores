`define MSG_OFFSET_EMPTY 0
`define MSG_OFFSET_STOPPED_TRAP 1
