@00000000
2B 3B 
24 23 30 30 3B 
24 53 30 30 23 42 33 3B
54 30 35
30 3A 30 30 30 30 3B
31 3A 31 31 31 31 3B
32 3A 32 32 32 32 3B
33 3A 33 33 33 33 3B
34 3A 34 34 34 34 3B
35 3A 35 35 35 35 3B
31 3A 30 30 30 30 3B
31 36 3A 30 30 30 30 3B
31 37 3A 30 30 30 30 3B

