@00000000
01 10 00 FF 9F A4 2E 00 01 20 00 00 1F 1C 01 30 
00 00 1F A4 2E 44 0E 23 C0 06 0D 24 00 00 82 04 
1A 00 00 00 10 16 01 20 00 00 FE ED 24 20 F0 00 
00 00 2E 22 2E 33 2E 44 03 00 00 00 19 B6 1A 00 
00 00 10 3E 01 30 00 00 00 01 22 20 F0 00 00 08 
0E 23 C7 FB 22 20 F0 00 00 0C 04 00 6D 6F 78 69 
65 00 91 18 01 30 00 00 1F 18 01 20 00 00 1F 18 
0E 32 C0 07 01 30 00 00 00 00 2E 44 0E 34 C0 01 
19 30 04 00 91 18 01 40 00 00 1F 18 01 20 00 00 
1F 18 29 42 01 30 00 00 00 02 2D 43 01 30 00 00 
00 1F 02 54 27 53 02 35 05 34 01 40 00 00 00 01 
2D 34 2E 55 0E 35 C0 06 01 40 00 00 00 00 0E 45 
C0 01 19 40 04 00 06 18 06 19 06 1A 91 18 1D 30 
00 00 1F 1C 2E 22 0E 32 C4 33 01 90 00 00 00 02 
01 80 00 00 1F 10 01 20 00 00 1F 0C 29 82 2D 89 
98 01 02 A2 08 20 00 00 1F 20 0E 28 E0 0E 82 01 
09 20 00 00 1F 20 28 29 02 3A 05 32 0A 23 19 20 
08 20 00 00 1F 20 0E 28 D3 F2 03 00 00 00 10 62 
01 30 00 00 00 00 2E 22 0E 32 C0 04 01 20 00 00 
1F 14 19 30 1B 20 00 00 00 01 1F 20 00 00 1F 1C 
02 E0 9E 0C 07 EA 07 E9 07 E8 04 00 91 18 04 00 
91 18 01 40 00 00 00 00 2E 22 0E 42 C0 07 01 30 
00 00 1F 24 01 20 00 00 1F 14 19 40 03 00 00 00 
10 84 04 00 91 18 04 00 01 30 F0 00 00 08 38 23 
00 02 11 22 01 40 00 00 00 01 0E 24 C0 05 38 23 
00 02 11 22 0E 24 C7 FB 20 20 00 00 00 23 39 32 
00 06 08 60 00 00 1F 9C 01 20 00 00 00 04 02 46 
2D 42 02 24 01 E0 00 00 00 0F 26 2E 01 40 00 00 
1E 1C 02 54 05 52 1C 55 01 20 00 00 1F 48 1E 25 
26 6E 05 46 1C 44 37 24 00 01 2E 44 37 24 00 02 
12 55 2E EE 0E 5E C0 12 02 42 01 60 00 00 00 01 
1A 00 00 00 11 F6 38 23 00 02 11 22 0E 26 C7 FB 
39 35 00 06 84 01 1C 54 0E 5E C7 F5 2E 22 09 20 
00 00 1F 9C 04 00 06 18 06 19 06 1A 06 1B 06 1C 
06 1D 91 18 02 92 99 01 2E DD 01 C0 00 00 10 44 
01 B0 00 00 00 46 01 A0 00 00 00 05 01 80 FF FF 
FF FF 1A 00 00 00 12 72 01 30 00 00 00 41 0E 43 
E0 20 92 30 12 22 01 50 00 00 00 09 0E 25 D4 15 
94 30 01 20 00 00 00 04 28 D2 05 D4 99 01 0E 98 
C0 14 19 C0 12 42 0E 4B E7 E7 92 61 12 22 0E 2A 
D4 04 94 57 1A 00 00 00 12 62 02 48 1A 00 00 00 
12 62 94 37 1A 00 00 00 12 62 02 2D 02 E0 9E 18 
07 ED 07 EC 07 EB 07 EA 07 E9 07 E8 04 00 06 18 
06 19 06 1A 06 1B 06 1C 06 1D 91 18 2E 88 01 D0 
00 00 10 44 01 C0 00 00 00 46 01 B0 00 00 00 05 
01 A0 00 00 00 41 01 90 00 00 00 09 19 D0 12 32 
0E 3C D4 12 0E 3A E0 18 92 30 12 22 0E 29 D4 18 
93 30 2E 22 0E 32 C8 14 01 20 00 00 00 04 28 82 
05 83 1A 00 00 00 12 DC 92 61 12 22 0E 2B D4 08 
93 57 1A 00 00 00 12 F2 93 37 1A 00 00 00 12 F2 
02 28 02 E0 9E 18 07 ED 07 EC 07 EB 07 EA 07 E9 
07 E8 04 00 06 18 06 19 06 1A 06 1B 06 1C 06 1D 
91 1C 01 80 F0 00 00 08 2E CC 01 90 00 00 00 01 
22 30 00 00 1F A0 11 23 0E 2C C1 19 24 C0 00 00 
1F A0 01 B0 00 00 10 44 19 B0 12 22 01 30 00 00 
00 63 0E 23 C0 F1 D4 76 01 30 00 00 00 4D 0E 23 
C4 03 1A 00 00 00 17 DE 01 30 00 00 00 50 0E 23 
C1 DC 01 30 00 00 00 3F 0E 23 C0 23 01 A0 00 00 
00 23 01 B0 00 00 10 44 19 B0 12 22 0E 2A C7 F9 
19 B0 19 B0 01 40 00 00 1E 3C 01 30 00 00 00 2B 
1A 00 00 00 13 C6 38 28 00 02 11 22 0E 29 C7 FB 
39 83 00 06 84 01 1C 34 0E 3C C7 F5 1A 00 00 00 
13 50 01 E0 00 00 10 44 19 E0 01 30 00 00 10 44 
19 30 01 40 00 00 10 44 19 40 01 40 00 00 1E 30 
01 30 00 00 00 2B 1A 00 00 00 14 0C 38 28 00 02 
11 22 0E 29 C7 FB 39 83 00 06 84 01 1C 34 0E 3C 
C7 F5 01 40 00 00 1E 38 01 30 00 00 00 53 1A 00 
00 00 14 34 38 28 00 02 11 22 0E 29 C7 FB 39 83 
00 06 08 20 00 00 1F 9C 05 23 09 20 00 00 1F 9C 
84 01 1C 34 0E 3C C7 EE 03 00 00 00 11 78 1A 00 
00 00 13 50 01 30 00 00 00 6D 0E 23 C1 05 01 30 
00 00 00 70 0E 23 C0 98 01 30 00 00 00 67 0E 23 
C7 8D 01 E0 00 00 10 44 19 E0 01 30 00 00 10 44 
19 30 01 40 00 00 10 44 19 40 01 40 00 00 1E 30 
01 30 00 00 00 2B 1A 00 00 00 14 AC 38 28 00 02 
11 22 0E 29 C7 FB 39 83 00 06 84 01 1C 34 0E 3C 
C7 F5 01 B0 00 00 1F 4C 01 D0 00 00 1F 3C 01 60 
00 00 1E 1C 01 A0 00 00 00 0F 01 70 FF FF FF FC 
0A 5B 01 40 00 00 1F 3C 01 20 00 00 00 1C 02 35 
2D 32 26 3A 02 E6 05 E3 1C 3E 1E 43 92 04 84 01 
0E 27 C7 F5 2E 22 37 D2 00 08 1C 3D 0E 3C C0 18 
01 40 00 00 1F 3C 1A 00 00 00 15 1C 38 28 00 02 
11 22 0E 29 C7 FB 39 83 00 06 08 20 00 00 1F 9C 
05 23 09 20 00 00 1F 9C 84 01 1C 34 0E 3C C7 EE 
8B 04 01 30 00 00 1F 94 0E B3 C7 CA 03 00 00 00 
11 78 1A 00 00 00 13 50 38 28 00 02 11 22 01 30 
00 00 00 01 0E 23 C0 05 38 28 00 02 11 22 0E 23 
C7 FB 20 20 00 00 00 2B 39 82 00 06 02 E0 9E 18 
07 ED 07 EC 07 EB 07 EA 07 E9 07 E8 04 00 01 A0 
00 00 00 24 01 40 00 00 10 44 19 40 12 22 0E 2A 
C7 F9 1A 00 00 00 13 62 03 00 00 00 12 AE 02 A2 
01 40 00 00 10 44 19 40 01 B0 00 00 10 44 19 B0 
01 40 00 00 1E 30 01 30 00 00 00 2B 1A 00 00 00 
15 D2 38 28 00 02 11 22 0E 29 C7 FB 39 83 00 06 
84 01 1C 34 0E 3C C7 F5 01 20 00 00 00 02 28 A2 
01 20 00 00 1F 4C 05 2A 0A A2 01 D0 00 00 1F 3C 
02 4D 01 20 00 00 00 1C 01 60 00 00 1E 1C 01 70 
00 00 00 0F 01 50 FF FF FF FC 02 3A 2D 32 26 37 
02 E6 05 E3 1C 3E 1E 43 92 04 84 01 0E 25 C7 F5 
2E 22 37 D2 00 08 1C 3D 0E 3C C3 0E 01 40 00 00 
1F 3C 1A 00 00 00 16 48 38 28 00 02 11 22 0E 29 
C7 FB 39 83 00 06 08 20 00 00 1F 9C 05 23 09 20 
00 00 1F 9C 84 01 1C 34 0E 3C C7 EE 03 00 00 00 
11 78 1A 00 00 00 13 50 01 A0 00 00 12 AE 19 A0 
02 B2 0D 02 FF E4 19 A0 02 A2 01 40 00 00 10 44 
19 40 01 E0 00 00 10 44 19 E0 01 50 00 00 1E 30 
01 40 00 00 00 2B 0C 30 FF E4 1A 00 00 00 16 B0 
38 28 00 02 11 22 0E 29 C7 FB 39 84 00 06 85 01 
1C 45 0E 4C C7 F5 05 AB 01 D0 00 00 00 04 01 60 
00 00 1E 1C 01 50 00 00 1F 48 01 B0 00 00 00 0F 
02 2A 29 23 0E 2C DE B8 02 73 87 01 1C 43 12 24 
2D 2D 02 36 05 32 1C 33 1E 53 02 2B 26 24 02 46 
05 42 1C 24 37 52 00 01 37 5C 00 02 12 33 0E 3C 
C0 18 01 40 00 00 1F 48 1A 00 00 00 17 1E 38 28 
00 02 11 22 0E 29 C7 FB 39 83 00 06 08 20 00 00 
1F 9C 05 23 09 20 00 00 1F 9C 84 01 1C 34 0E 3C 
C7 EE 02 37 1A 00 00 00 16 E0 01 B0 00 00 12 AE 
19 B0 02 A2 19 B0 01 30 00 00 00 02 02 4A 28 43 
01 30 00 00 1F 4C 05 34 0B 32 01 B0 00 00 10 44 
19 B0 19 B0 01 40 00 00 1E 30 01 30 00 00 00 2B 
1A 00 00 00 17 86 38 28 00 02 11 22 0E 29 C7 FB 
39 83 00 06 84 01 1C 34 0E 3C C7 F5 01 40 00 00 
1E 34 01 30 00 00 00 4F 1A 00 00 00 17 AE 38 28 
00 02 11 22 0E 29 C7 FB 39 83 00 06 08 20 00 00 
1F 9C 05 23 09 20 00 00 1F 9C 84 01 1C 34 0E 3C 
C7 EE 03 00 00 00 11 78 1A 00 00 00 13 50 01 A0 
00 00 12 AE 19 A0 02 B2 19 A0 0E 2C DC 0D 02 A2 
05 AB 01 D0 00 00 12 16 01 20 00 00 00 02 19 D0 
1E B2 8B 01 0E BA C7 F8 01 40 00 00 1E 30 01 30 
00 00 00 2B 1A 00 00 00 18 1A 38 28 00 02 11 22 
0E 29 C7 FB 39 83 00 06 84 01 1C 34 0E 3C C7 F5 
01 40 00 00 1E 34 01 30 00 00 00 4F 1A 00 00 00 
18 42 38 28 00 02 11 22 0E 29 C7 FB 39 83 00 06 
08 20 00 00 1F 9C 05 23 09 20 00 00 1F 9C 84 01 
1C 34 0E 3C C7 EE 03 00 00 00 11 78 1A 00 00 00 
13 50 06 18 06 19 06 1A 06 1B 06 1C 91 1C 01 40 
00 00 00 05 0E 34 D4 26 01 40 00 00 00 01 02 54 
28 53 02 35 01 50 00 00 00 1B 02 63 26 65 2E 55 
0E 65 C4 21 01 50 00 00 00 20 02 83 26 85 0E 86 
C4 20 01 40 00 00 00 04 26 34 0E 38 C0 0B 24 80 
F0 00 00 10 02 E0 9E 14 07 EC 07 EB 07 EA 07 E9 
07 E8 04 00 20 20 FF FF FF FF 24 20 F0 00 00 00 
1A 00 00 00 18 E0 24 50 F0 00 00 00 1A 00 00 00 
18 EC 02 B0 01 30 F0 00 00 08 38 53 00 02 11 55 
0E 54 C0 05 38 53 00 02 11 55 0E 54 C7 FB 20 40 
00 00 00 24 39 34 00 06 01 50 00 00 1E 38 01 40 
00 00 00 53 01 70 00 00 00 01 2E 88 1A 00 00 00 
19 32 38 63 00 02 11 66 0E 67 C7 FB 39 34 00 06 
08 60 00 00 1F 9C 05 64 09 60 00 00 1F 9C 85 01 
1C 45 0E 48 C7 EE 0D 02 FF E8 03 00 00 00 11 78 
02 AB 8A 0C 01 80 00 00 1F 54 02 C8 8C 38 02 38 
02 4A 0C 20 FF E8 0A 54 0B 35 84 04 83 04 0E 3C 
C7 FA 0A 3B 01 90 00 00 1F 4C 0D 93 00 04 0A 3B 
0A 33 0B 93 92 02 0D 92 00 40 03 00 00 00 13 34 
0A 28 0B A2 88 04 8A 04 0E 8C C7 FA 0C 29 00 40 
1A 00 00 00 18 C4 06 18 06 19 06 1A 06 1B 06 1C 
06 1D 91 30 01 80 F0 00 00 08 20 20 00 00 00 58 
39 82 00 06 20 20 00 00 00 59 39 82 00 06 20 20 
00 00 00 5A 39 82 00 06 01 20 00 00 1D 70 B2 01 
01 30 00 00 00 01 B3 00 2E 22 09 20 00 00 1F 9C 
01 60 00 00 1E 44 01 50 00 00 00 4D 02 42 1A 00 
00 00 1A 14 38 28 00 02 11 22 0E 23 C7 FB 39 85 
00 06 86 01 1C 56 0E 54 C7 F5 01 50 00 00 1E 64 
01 40 00 00 00 43 01 30 00 00 00 01 2E 66 1A 00 
00 00 1A 44 38 28 00 02 11 22 0E 23 C7 FB 39 84 
00 06 85 01 1C 45 0E 46 C7 F5 01 50 00 00 1E DC 
01 40 00 00 00 0A 01 30 00 00 00 01 2E 66 1A 00 
00 00 1A 74 38 28 00 02 11 22 0E 23 C7 FB 39 84 
00 06 85 01 1C 45 0E 46 C7 F5 01 50 00 00 1E A0 
01 40 00 00 00 57 01 30 00 00 00 01 2E 66 1A 00 
00 00 1A A4 38 28 00 02 11 22 0E 23 C7 FB 39 84 
00 06 85 01 1C 45 0E 46 C7 F5 20 20 00 00 00 01 
24 20 00 00 1F A0 01 B0 00 00 10 44 01 A0 00 00 
00 24 01 90 00 00 00 53 1A 00 00 00 1A E2 0E 29 
C0 1B 19 B0 12 22 0E 2A C7 FA 20 20 FF FF DE B2 
24 20 F0 00 00 00 01 80 00 00 1F 4C 02 28 02 48 
84 50 2E 33 0B 23 82 04 0E 42 C7 FC 03 00 00 00 
13 34 0C 88 00 40 25 80 20 A0 00 00 00 01 01 C0 
00 00 12 16 22 30 00 00 1F A0 11 23 2E 44 0E 24 
C0 5C 2E 44 24 40 00 00 1F A0 19 B0 12 D2 02 3D 
02 2D 92 30 13 22 01 40 00 00 00 09 0E 24 D5 03 
01 20 00 00 00 02 0D 03 FF E0 19 C0 02 92 24 A0 
F0 00 00 00 01 20 00 00 00 33 0E D2 0C 30 FF E0 
C0 67 E4 4C 01 20 00 00 00 37 0E D2 C0 D8 01 20 
00 00 00 39 0E D2 C4 C6 21 38 11 33 2E 22 0E 32 
C0 08 38 38 00 04 39 03 FF E6 21 38 11 33 0E 32 
C7 F8 01 30 00 00 1E E0 01 20 00 00 00 4A 01 50 
00 00 00 01 2E 66 1A 00 00 00 1B BC 38 48 00 02 
11 44 0E 45 C7 FB 39 82 00 06 83 01 1C 23 0E 26 
C7 F5 20 20 00 00 30 00 24 20 F0 00 00 00 1A 00 
30 00 00 00 1A 00 00 00 1B E4 19 B0 12 22 01 30 
00 00 00 53 0E 23 C3 A1 19 B0 12 22 01 30 00 00 
00 53 0E 23 C7 F2 1A 00 00 00 1B 3A 01 20 00 00 
00 30 0E D2 C4 7F 05 99 02 D9 9D 01 8A 01 13 99 
2E 33 0E 93 C3 7F 01 90 FF FF FF FF 19 B0 02 2D 
92 01 02 D2 11 22 0E 29 C7 F9 1A 00 00 00 1B 24 
01 20 00 00 00 08 19 C0 02 32 02 49 94 04 02 D4 
11 54 01 20 00 00 00 04 0E 52 DC 36 02 D9 9D 09 
13 DD 01 20 00 00 00 02 27 D2 13 9D 02 59 28 52 
85 04 05 53 02 63 01 70 00 00 00 08 02 27 0D 03 
FF E0 0D 04 FF D0 0D 05 FF D8 0D 06 FF D4 0D 07 
FF DC 19 C0 0C 60 FF D4 0B 62 86 04 0C 50 FF D8 
0E 56 0C 30 FF E0 0C 40 FF D0 0C 70 FF DC C7 E6 
02 29 82 01 01 50 00 00 00 02 28 25 05 32 28 D5 
02 24 29 2D 92 04 02 D2 11 2D 01 40 00 00 00 02 
0E 24 DC 0D 01 20 00 00 00 04 0D 03 FF E0 19 C0 
0C 30 FF E0 23 32 83 02 02 2D 92 02 11 22 01 40 
00 00 00 02 0E 24 C4 06 0D 03 FF E0 19 C0 0C 30 
FF E0 1E 32 01 20 00 00 00 02 19 C0 8A 01 1A 00 
00 00 1B 24 01 20 00 00 00 08 02 43 28 42 02 24 
05 2A 24 20 F0 00 00 00 1A 00 00 00 1D 28 05 99 
02 A9 9A 01 13 99 2E 22 0E 92 C3 26 01 90 FF FF 
FF FF 19 B0 02 2A 92 01 02 A2 11 22 0E 29 C7 F9 
1A 00 00 00 1B 88 01 20 00 00 00 08 02 43 28 42 
02 24 05 2A 24 20 F0 00 00 00 1A 00 00 00 1D 6A 
91 0C 0B 10 02 01 06 1F 06 1E 06 1D 06 1C 06 1B 
06 1A 06 19 06 18 06 17 06 16 06 15 06 14 06 13 
06 12 A2 05 A3 02 A4 03 03 00 00 00 18 72 0D 02 
00 04 01 60 00 00 00 01 A5 00 2B 56 B5 00 02 20 
92 38 02 12 07 12 07 13 07 14 07 15 07 16 07 17 
07 18 07 19 07 1A 07 1B 07 1C 07 1D 07 1E 07 1F 
04 00 06 18 06 19 91 18 01 80 00 00 1F 08 0C 28 
FF FC 01 90 FF FF FF FF 0E 29 C0 06 98 04 19 20 
98 04 0A 28 0E 29 C7 FB 02 E0 9E 08 07 E9 07 E8 
04 00 91 18 04 00 03 00 00 00 11 50 03 00 00 00 
1D D2 04 00 03 00 00 00 10 C6 04 00 
@00000E1C
30 31 32 33 34 35 36 37 38 39 41 42 43 44 45 46 
00 00 00 00 2B 24 00 00 4F 4B 00 00 53 30 35 00 
2B 24 23 30 30 00 00 00 4D 4F 58 49 45 20 4F 6E 
2D 43 68 69 70 20 42 6F 6F 74 6C 6F 61 64 65 72 
20 76 32 2E 30 0A 0D 00 43 6F 70 79 72 69 67 68 
74 20 28 63 29 20 32 30 31 33 20 41 6E 74 68 6F 
6E 79 20 47 72 65 65 6E 20 3C 67 72 65 65 6E 40 
6D 6F 78 69 65 6C 6F 67 69 63 2E 63 6F 6D 3E 0A 
0D 00 00 00 57 61 69 74 69 6E 67 20 66 6F 72 20 
61 6E 20 53 2D 52 65 63 6F 72 64 20 44 6F 77 6E 
6C 6F 61 64 20 6F 72 20 52 65 6D 6F 74 65 20 47 
44 42 20 43 6F 6E 6E 65 63 74 69 6F 6E 2E 2E 2E 
0A 0D 00 00 4A 75 6D 70 69 6E 67 20 74 6F 20 63 
6F 64 65 20 61 74 20 30 78 33 30 30 30 30 30 30 
30 2E 0A 0D 00 00 00 00 FF FF FF FF 00 00 00 00 
FF FF FF FF 00 00 00 00 00 00 00 00 
@00000F18
00 00 00 00 
